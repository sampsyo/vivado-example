/* verilator lint_off PINMISSING */
/* verilator lint_off WIDTH */
module std_mem_d2
  #(parameter width = 32,
    parameter d0_size = 16,
    parameter d1_size = 16,
    parameter d0_idx_size = 4,
    parameter d1_idx_size = 4)
   (input logic [d0_idx_size-1:0] addr0,
    input logic [d1_idx_size-1:0] addr1,
    input logic [width-1:0]   write_data,
    input logic               write_en,
    input logic               clk,
    output logic [width-1:0]  read_data,
    output logic done);

  logic [width-1:0]  mem[d0_size-1:0][d1_size-1:0];

  assign read_data = mem[addr0][addr1];
  always_ff @(posedge clk) begin
    if (write_en) begin
      mem[addr0][addr1] <= write_data;
      done <= 1'd1;
    end else
      done <= 1'd0;
  end
endmodule

module std_add
  #(parameter width = 32)
  (input  logic [width-1:0] left,
    input  logic [width-1:0] right,
    output logic [width-1:0] out);
  assign out = left + right;
endmodule

module std_reg
  #(parameter width = 32)
   (input wire [width-1:0] in,
    input wire write_en,
    input wire clk,
    // output
    output logic [width - 1:0] out,
    output logic done);

  always_ff @(posedge clk) begin
    if (write_en) begin
      out <= in;
      done <= 1'd1;
    end else
      done <= 1'd0;
  end
endmodule

module std_const
  #(parameter width = 32,
    parameter value = 0)
   (input logic                valid,
    output logic               ready,
    output logic [width - 1:0] out,
    output logic               out_read_out);
  assign out = value;
  assign ready = valid;
  assign out_read_out = valid;
endmodule

module std_le
  #(parameter width = 32)
  (input logic [width-1:0] left,
   input logic [width-1:0] right,
   output logic            out);
  assign out = left <= right;
endmodule

module std_mult
  #(parameter width = 32)
  (input logic  [width-1:0] left,
    input logic  [width-1:0] right,
    output logic [width-1:0] out);
  assign out = left * right;
endmodule

module std_mem_d1
  #(parameter width = 32,
    parameter size = 16,
    parameter idx_size = 4)
   (input logic [idx_size-1:0] addr0,
    input logic [width-1:0]   write_data,
    input logic               write_en,
    input logic               clk,
    output logic [width-1:0]  read_data,
    output logic done);

  logic [width-1:0]  mem[size-1:0];

  assign read_data = mem[addr0];
  always_ff @(posedge clk) begin
    if (write_en) begin
      mem[addr0] <= write_data;
      done <= 1'd1;
    end else
      done <= 1'd0;
  end
endmodule

// Component Signature
module main (
      input wire clk,
      input wire go,
      output wire done
  );
  
  // Structure wire declarations
  wire [3:0] A_addr0;
  wire [3:0] A_addr1;
  wire [31:0] A_write_data;
  wire A_write_en;
  wire A_clk;
  wire [31:0] A_read_data;
  wire A_done;
  wire [3:0] add0_left;
  wire [3:0] add0_right;
  wire [3:0] add0_out;
  wire [31:0] add1_left;
  wire [31:0] add1_right;
  wire [31:0] add1_out;
  wire [3:0] add2_left;
  wire [3:0] add2_right;
  wire [3:0] add2_out;
  wire [31:0] add3_left;
  wire [31:0] add3_right;
  wire [31:0] add3_out;
  wire [3:0] add4_left;
  wire [3:0] add4_right;
  wire [3:0] add4_out;
  wire [3:0] add5_left;
  wire [3:0] add5_right;
  wire [3:0] add5_out;
  wire const0_valid;
  wire [3:0] const0_out;
  wire const0_out_read_out;
  wire const0_ready;
  wire const1_valid;
  wire [3:0] const1_out;
  wire const1_out_read_out;
  wire const1_ready;
  wire const10_valid;
  wire [3:0] const10_out;
  wire const10_out_read_out;
  wire const10_ready;
  wire const11_valid;
  wire [3:0] const11_out;
  wire const11_out_read_out;
  wire const11_ready;
  wire const12_valid;
  wire [3:0] const12_out;
  wire const12_out_read_out;
  wire const12_ready;
  wire const13_valid;
  wire [3:0] const13_out;
  wire const13_out_read_out;
  wire const13_ready;
  wire const2_valid;
  wire [31:0] const2_out;
  wire const2_out_read_out;
  wire const2_ready;
  wire const3_valid;
  wire [3:0] const3_out;
  wire const3_out_read_out;
  wire const3_ready;
  wire const4_valid;
  wire [3:0] const4_out;
  wire const4_out_read_out;
  wire const4_ready;
  wire const5_valid;
  wire [3:0] const5_out;
  wire const5_out_read_out;
  wire const5_ready;
  wire const6_valid;
  wire [31:0] const6_out;
  wire const6_out_read_out;
  wire const6_ready;
  wire const7_valid;
  wire [3:0] const7_out;
  wire const7_out_read_out;
  wire const7_ready;
  wire const8_valid;
  wire [3:0] const8_out;
  wire const8_out_read_out;
  wire const8_ready;
  wire const9_valid;
  wire [3:0] const9_out;
  wire const9_out_read_out;
  wire const9_ready;
  wire [3:0] i0_in;
  wire i0_write_en;
  wire i0_clk;
  wire [3:0] i0_out;
  wire i0_done;
  wire [3:0] i1_in;
  wire i1_write_en;
  wire i1_clk;
  wire [3:0] i1_out;
  wire i1_done;
  wire [3:0] j0_in;
  wire j0_write_en;
  wire j0_clk;
  wire [3:0] j0_out;
  wire j0_done;
  wire [3:0] j1_in;
  wire j1_write_en;
  wire j1_clk;
  wire [3:0] j1_out;
  wire j1_done;
  wire [3:0] le0_left;
  wire [3:0] le0_right;
  wire le0_out;
  wire [3:0] le1_left;
  wire [3:0] le1_right;
  wire le1_out;
  wire [3:0] le2_left;
  wire [3:0] le2_right;
  wire le2_out;
  wire [3:0] le3_left;
  wire [3:0] le3_right;
  wire le3_out;
  wire [31:0] mult0_left;
  wire [31:0] mult0_right;
  wire [31:0] mult0_out;
  wire [31:0] mult1_left;
  wire [31:0] mult1_right;
  wire [31:0] mult1_out;
  wire [31:0] t0_in;
  wire t0_write_en;
  wire t0_clk;
  wire [31:0] t0_out;
  wire t0_done;
  wire [3:0] tmp_addr0;
  wire [31:0] tmp_write_data;
  wire tmp_write_en;
  wire tmp_clk;
  wire [31:0] tmp_read_data;
  wire tmp_done;
  wire [3:0] x_addr0;
  wire [31:0] x_write_data;
  wire x_write_en;
  wire x_clk;
  wire [31:0] x_read_data;
  wire x_done;
  wire [3:0] y_addr0;
  wire [31:0] y_write_data;
  wire y_write_en;
  wire y_clk;
  wire [31:0] y_read_data;
  wire y_done;
  wire [31:0] y00_in;
  wire y00_write_en;
  wire y00_clk;
  wire [31:0] y00_out;
  wire y00_done;
  wire [31:0] fsm0_in;
  wire fsm0_write_en;
  wire fsm0_clk;
  wire [31:0] fsm0_out;
  wire fsm0_done;
  wire [31:0] incr0_left;
  wire [31:0] incr0_right;
  wire [31:0] incr0_out;
  wire [31:0] fsm1_in;
  wire fsm1_write_en;
  wire fsm1_clk;
  wire [31:0] fsm1_out;
  wire fsm1_done;
  wire cond_stored0_in;
  wire cond_stored0_write_en;
  wire cond_stored0_clk;
  wire cond_stored0_out;
  wire cond_stored0_done;
  wire [31:0] incr1_left;
  wire [31:0] incr1_right;
  wire [31:0] incr1_out;
  wire [31:0] fsm2_in;
  wire fsm2_write_en;
  wire fsm2_clk;
  wire [31:0] fsm2_out;
  wire fsm2_done;
  wire [31:0] incr2_left;
  wire [31:0] incr2_right;
  wire [31:0] incr2_out;
  wire [31:0] fsm3_in;
  wire fsm3_write_en;
  wire fsm3_clk;
  wire [31:0] fsm3_out;
  wire fsm3_done;
  wire cond_stored1_in;
  wire cond_stored1_write_en;
  wire cond_stored1_clk;
  wire cond_stored1_out;
  wire cond_stored1_done;
  wire [31:0] incr3_left;
  wire [31:0] incr3_right;
  wire [31:0] incr3_out;
  wire [31:0] fsm4_in;
  wire fsm4_write_en;
  wire fsm4_clk;
  wire [31:0] fsm4_out;
  wire fsm4_done;
  wire [31:0] incr4_left;
  wire [31:0] incr4_right;
  wire [31:0] incr4_out;
  wire [31:0] fsm5_in;
  wire fsm5_write_en;
  wire fsm5_clk;
  wire [31:0] fsm5_out;
  wire fsm5_done;
  wire cond_stored2_in;
  wire cond_stored2_write_en;
  wire cond_stored2_clk;
  wire cond_stored2_out;
  wire cond_stored2_done;
  wire [31:0] incr5_left;
  wire [31:0] incr5_right;
  wire [31:0] incr5_out;
  wire [31:0] fsm6_in;
  wire fsm6_write_en;
  wire fsm6_clk;
  wire [31:0] fsm6_out;
  wire fsm6_done;
  wire cond_computed0_in;
  wire cond_computed0_write_en;
  wire cond_computed0_clk;
  wire cond_computed0_out;
  wire cond_computed0_done;
  wire cond_stored3_in;
  wire cond_stored3_write_en;
  wire cond_stored3_clk;
  wire cond_stored3_out;
  wire cond_stored3_done;
  wire done_reg0_in;
  wire done_reg0_write_en;
  wire done_reg0_clk;
  wire done_reg0_out;
  wire done_reg0_done;
  wire [31:0] fsm7_in;
  wire fsm7_write_en;
  wire fsm7_clk;
  wire [31:0] fsm7_out;
  wire fsm7_done;
  
  // Subcomponent Instances
  std_mem_d2 #(32, 8, 8, 4, 4) A (
      .addr0(A_addr0),
      .addr1(A_addr1),
      .clk(clk),
      .read_data(A_read_data),
      .done(A_done)
  );
  
  std_add #(4) add0 (
      .left(add0_left),
      .right(add0_right),
      .out(add0_out)
  );
  
  std_add #(32) add1 (
      .left(add1_left),
      .right(add1_right),
      .out(add1_out)
  );
  
  std_add #(4) add2 (
      .left(add2_left),
      .right(add2_right),
      .out(add2_out)
  );
  
  std_add #(32) add3 (
      .left(add3_left),
      .right(add3_right),
      .out(add3_out)
  );
  
  std_add #(4) add4 (
      .left(add4_left),
      .right(add4_right),
      .out(add4_out)
  );
  
  std_add #(4) add5 (
      .left(add5_left),
      .right(add5_right),
      .out(add5_out)
  );
  
  std_const #(4, 0) const0 (
      .out(const0_out),
      .out_read_out(const0_out_read_out),
      .ready(const0_ready)
  );
  
  std_const #(4, 7) const1 (
      .out(const1_out),
      .out_read_out(const1_out_read_out),
      .ready(const1_ready)
  );
  
  std_const #(4, 0) const10 (
      .out(const10_out),
      .out_read_out(const10_out_read_out),
      .ready(const10_ready)
  );
  
  std_const #(4, 7) const11 (
      .out(const11_out),
      .out_read_out(const11_out_read_out),
      .ready(const11_ready)
  );
  
  std_const #(4, 1) const12 (
      .out(const12_out),
      .out_read_out(const12_out_read_out),
      .ready(const12_ready)
  );
  
  std_const #(4, 1) const13 (
      .out(const13_out),
      .out_read_out(const13_out_read_out),
      .ready(const13_ready)
  );
  
  std_const #(32, 0) const2 (
      .out(const2_out),
      .out_read_out(const2_out_read_out),
      .ready(const2_ready)
  );
  
  std_const #(4, 1) const3 (
      .out(const3_out),
      .out_read_out(const3_out_read_out),
      .ready(const3_ready)
  );
  
  std_const #(4, 0) const4 (
      .out(const4_out),
      .out_read_out(const4_out_read_out),
      .ready(const4_ready)
  );
  
  std_const #(4, 7) const5 (
      .out(const5_out),
      .out_read_out(const5_out_read_out),
      .ready(const5_ready)
  );
  
  std_const #(32, 0) const6 (
      .out(const6_out),
      .out_read_out(const6_out_read_out),
      .ready(const6_ready)
  );
  
  std_const #(4, 0) const7 (
      .out(const7_out),
      .out_read_out(const7_out_read_out),
      .ready(const7_ready)
  );
  
  std_const #(4, 7) const8 (
      .out(const8_out),
      .out_read_out(const8_out_read_out),
      .ready(const8_ready)
  );
  
  std_const #(4, 1) const9 (
      .out(const9_out),
      .out_read_out(const9_out_read_out),
      .ready(const9_ready)
  );
  
  std_reg #(4) i0 (
      .in(i0_in),
      .write_en(i0_write_en),
      .clk(clk),
      .out(i0_out),
      .done(i0_done)
  );
  
  std_reg #(4) i1 (
      .in(i1_in),
      .write_en(i1_write_en),
      .clk(clk),
      .out(i1_out),
      .done(i1_done)
  );
  
  std_reg #(4) j0 (
      .in(j0_in),
      .write_en(j0_write_en),
      .clk(clk),
      .out(j0_out),
      .done(j0_done)
  );
  
  std_reg #(4) j1 (
      .in(j1_in),
      .write_en(j1_write_en),
      .clk(clk),
      .out(j1_out),
      .done(j1_done)
  );
  
  std_le #(4) le0 (
      .left(le0_left),
      .right(le0_right),
      .out(le0_out)
  );
  
  std_le #(4) le1 (
      .left(le1_left),
      .right(le1_right),
      .out(le1_out)
  );
  
  std_le #(4) le2 (
      .left(le2_left),
      .right(le2_right),
      .out(le2_out)
  );
  
  std_le #(4) le3 (
      .left(le3_left),
      .right(le3_right),
      .out(le3_out)
  );
  
  std_mult #(32) mult0 (
      .left(mult0_left),
      .right(mult0_right),
      .out(mult0_out)
  );
  
  std_mult #(32) mult1 (
      .left(mult1_left),
      .right(mult1_right),
      .out(mult1_out)
  );
  
  std_reg #(32) t0 (
      .in(t0_in),
      .write_en(t0_write_en),
      .clk(clk),
      .out(t0_out),
      .done(t0_done)
  );
  
  std_mem_d1 #(32, 8, 4) tmp (
      .addr0(tmp_addr0),
      .write_data(tmp_write_data),
      .write_en(tmp_write_en),
      .clk(clk),
      .read_data(tmp_read_data),
      .done(tmp_done)
  );
  
  std_mem_d1 #(32, 8, 4) x (
      .addr0(x_addr0),
      .clk(clk),
      .read_data(x_read_data),
      .done(x_done)
  );
  
  std_mem_d1 #(32, 8, 4) y (
      .addr0(y_addr0),
      .write_data(y_write_data),
      .write_en(y_write_en),
      .clk(clk),
      .read_data(y_read_data),
      .done(y_done)
  );
  
  std_reg #(32) y00 (
      .in(y00_in),
      .write_en(y00_write_en),
      .clk(clk),
      .out(y00_out),
      .done(y00_done)
  );
  
  std_reg #(32) fsm0 (
      .in(fsm0_in),
      .write_en(fsm0_write_en),
      .clk(clk),
      .out(fsm0_out),
      .done(fsm0_done)
  );
  
  std_add #(32) incr0 (
      .left(incr0_left),
      .right(incr0_right),
      .out(incr0_out)
  );
  
  std_reg #(32) fsm1 (
      .in(fsm1_in),
      .write_en(fsm1_write_en),
      .clk(clk),
      .out(fsm1_out),
      .done(fsm1_done)
  );
  
  std_reg #(1) cond_stored0 (
      .in(cond_stored0_in),
      .write_en(cond_stored0_write_en),
      .clk(clk),
      .out(cond_stored0_out),
      .done(cond_stored0_done)
  );
  
  std_add #(32) incr1 (
      .left(incr1_left),
      .right(incr1_right),
      .out(incr1_out)
  );
  
  std_reg #(32) fsm2 (
      .in(fsm2_in),
      .write_en(fsm2_write_en),
      .clk(clk),
      .out(fsm2_out),
      .done(fsm2_done)
  );
  
  std_add #(32) incr2 (
      .left(incr2_left),
      .right(incr2_right),
      .out(incr2_out)
  );
  
  std_reg #(32) fsm3 (
      .in(fsm3_in),
      .write_en(fsm3_write_en),
      .clk(clk),
      .out(fsm3_out),
      .done(fsm3_done)
  );
  
  std_reg #(1) cond_stored1 (
      .in(cond_stored1_in),
      .write_en(cond_stored1_write_en),
      .clk(clk),
      .out(cond_stored1_out),
      .done(cond_stored1_done)
  );
  
  std_add #(32) incr3 (
      .left(incr3_left),
      .right(incr3_right),
      .out(incr3_out)
  );
  
  std_reg #(32) fsm4 (
      .in(fsm4_in),
      .write_en(fsm4_write_en),
      .clk(clk),
      .out(fsm4_out),
      .done(fsm4_done)
  );
  
  std_add #(32) incr4 (
      .left(incr4_left),
      .right(incr4_right),
      .out(incr4_out)
  );
  
  std_reg #(32) fsm5 (
      .in(fsm5_in),
      .write_en(fsm5_write_en),
      .clk(clk),
      .out(fsm5_out),
      .done(fsm5_done)
  );
  
  std_reg #(1) cond_stored2 (
      .in(cond_stored2_in),
      .write_en(cond_stored2_write_en),
      .clk(clk),
      .out(cond_stored2_out),
      .done(cond_stored2_done)
  );
  
  std_add #(32) incr5 (
      .left(incr5_left),
      .right(incr5_right),
      .out(incr5_out)
  );
  
  std_reg #(32) fsm6 (
      .in(fsm6_in),
      .write_en(fsm6_write_en),
      .clk(clk),
      .out(fsm6_out),
      .done(fsm6_done)
  );
  
  std_reg #(1) cond_computed0 (
      .in(cond_computed0_in),
      .write_en(cond_computed0_write_en),
      .clk(clk),
      .out(cond_computed0_out),
      .done(cond_computed0_done)
  );
  
  std_reg #(1) cond_stored3 (
      .in(cond_stored3_in),
      .write_en(cond_stored3_write_en),
      .clk(clk),
      .out(cond_stored3_out),
      .done(cond_stored3_done)
  );
  
  std_reg #(1) done_reg0 (
      .in(done_reg0_in),
      .write_en(done_reg0_write_en),
      .clk(clk),
      .out(done_reg0_out),
      .done(done_reg0_done)
  );
  
  std_reg #(32) fsm7 (
      .in(fsm7_in),
      .write_en(fsm7_write_en),
      .clk(clk),
      .out(fsm7_out),
      .done(fsm7_done)
  );
  
  
  // Input / output connections
  assign done = (fsm7_out == 32'd4) ? 1'd1 : '0;
  assign A_addr0 = (fsm2_out == 32'd1 & cond_stored1_out & fsm3_out >= 32'd1 & fsm3_out < 32'd4 & fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go | fsm4_out == 32'd1 & cond_stored2_out & fsm5_out >= 32'd1 & fsm5_out < 32'd4 & fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? i1_out : '0;
  assign A_addr1 = (fsm4_out == 32'd1 & cond_stored2_out & fsm5_out >= 32'd1 & fsm5_out < 32'd4 & fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? j1_out : (fsm2_out == 32'd1 & cond_stored1_out & fsm3_out >= 32'd1 & fsm3_out < 32'd4 & fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? j0_out : '0;
  assign add0_left = (fsm0_out == 32'd1 & cond_stored0_out & fsm1_out >= 32'd1 & fsm1_out < 32'd3 & fsm7_out == 32'd1 & !(fsm1_out == 32'd1 & !cond_stored0_out) & go) ? i0_out : '0;
  assign add0_right = (fsm0_out == 32'd1 & cond_stored0_out & fsm1_out >= 32'd1 & fsm1_out < 32'd3 & fsm7_out == 32'd1 & !(fsm1_out == 32'd1 & !cond_stored0_out) & go) ? const3_out : '0;
  assign add1_left = (fsm2_out == 32'd1 & cond_stored1_out & fsm3_out >= 32'd1 & fsm3_out < 32'd4 & fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? t0_out : '0;
  assign add1_right = (fsm2_out == 32'd1 & cond_stored1_out & fsm3_out >= 32'd1 & fsm3_out < 32'd4 & fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? mult0_out : '0;
  assign add2_left = (fsm2_out == 32'd2 & cond_stored1_out & fsm3_out >= 32'd1 & fsm3_out < 32'd4 & fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? j0_out : '0;
  assign add2_right = (fsm2_out == 32'd2 & cond_stored1_out & fsm3_out >= 32'd1 & fsm3_out < 32'd4 & fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? const9_out : '0;
  assign add3_left = (fsm4_out == 32'd1 & cond_stored2_out & fsm5_out >= 32'd1 & fsm5_out < 32'd4 & fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? y00_out : '0;
  assign add3_right = (fsm4_out == 32'd1 & cond_stored2_out & fsm5_out >= 32'd1 & fsm5_out < 32'd4 & fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? mult1_out : '0;
  assign add4_left = (fsm4_out == 32'd2 & cond_stored2_out & fsm5_out >= 32'd1 & fsm5_out < 32'd4 & fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? j1_out : '0;
  assign add4_right = (fsm4_out == 32'd2 & cond_stored2_out & fsm5_out >= 32'd1 & fsm5_out < 32'd4 & fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? const12_out : '0;
  assign add5_left = (fsm6_out == 32'd5 & !i1_done & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? i1_out : '0;
  assign add5_right = (fsm6_out == 32'd5 & !i1_done & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? const13_out : '0;
  assign i0_in = (fsm7_out == 32'd0 & !i0_done & go) ? const0_out : (fsm0_out == 32'd1 & cond_stored0_out & fsm1_out >= 32'd1 & fsm1_out < 32'd3 & fsm7_out == 32'd1 & !(fsm1_out == 32'd1 & !cond_stored0_out) & go) ? add0_out : '0;
  assign i0_write_en = (fsm7_out == 32'd0 & !i0_done & go | fsm0_out == 32'd1 & cond_stored0_out & fsm1_out >= 32'd1 & fsm1_out < 32'd3 & fsm7_out == 32'd1 & !(fsm1_out == 32'd1 & !cond_stored0_out) & go) ? 1'd1 : '0;
  assign i1_in = (fsm7_out == 32'd2 & !i1_done & go) ? const4_out : (fsm6_out == 32'd5 & !i1_done & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? add5_out : '0;
  assign i1_write_en = (fsm7_out == 32'd2 & !i1_done & go | fsm6_out == 32'd5 & !i1_done & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? 1'd1 : '0;
  assign j0_in = (fsm6_out == 32'd1 & !j0_done & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? const7_out : (fsm2_out == 32'd2 & cond_stored1_out & fsm3_out >= 32'd1 & fsm3_out < 32'd4 & fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? add2_out : '0;
  assign j0_write_en = (fsm6_out == 32'd1 & !j0_done & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go | fsm2_out == 32'd2 & cond_stored1_out & fsm3_out >= 32'd1 & fsm3_out < 32'd4 & fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? 1'd1 : '0;
  assign j1_in = (fsm6_out == 32'd3 & !j1_done & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? const10_out : (fsm4_out == 32'd2 & cond_stored2_out & fsm5_out >= 32'd1 & fsm5_out < 32'd4 & fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? add4_out : '0;
  assign j1_write_en = (fsm6_out == 32'd3 & !j1_done & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go | fsm4_out == 32'd2 & cond_stored2_out & fsm5_out >= 32'd1 & fsm5_out < 32'd4 & fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? 1'd1 : '0;
  assign le0_left = (fsm1_out < 32'd1 & fsm7_out == 32'd1 & !(fsm1_out == 32'd1 & !cond_stored0_out) & go) ? i0_out : '0;
  assign le0_right = (fsm1_out < 32'd1 & fsm7_out == 32'd1 & !(fsm1_out == 32'd1 & !cond_stored0_out) & go) ? const1_out : '0;
  assign le1_left = (!cond_computed0_out & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? i1_out : '0;
  assign le1_right = (!cond_computed0_out & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? const5_out : '0;
  assign le2_left = (fsm3_out < 32'd1 & fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? j0_out : '0;
  assign le2_right = (fsm3_out < 32'd1 & fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? const8_out : '0;
  assign le3_left = (fsm5_out < 32'd1 & fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? j1_out : '0;
  assign le3_right = (fsm5_out < 32'd1 & fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? const11_out : '0;
  assign mult0_left = (fsm2_out == 32'd1 & cond_stored1_out & fsm3_out >= 32'd1 & fsm3_out < 32'd4 & fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? A_read_data : '0;
  assign mult0_right = (fsm2_out == 32'd1 & cond_stored1_out & fsm3_out >= 32'd1 & fsm3_out < 32'd4 & fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? x_read_data : '0;
  assign mult1_left = (fsm4_out == 32'd1 & cond_stored2_out & fsm5_out >= 32'd1 & fsm5_out < 32'd4 & fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? A_read_data : '0;
  assign mult1_right = (fsm4_out == 32'd1 & cond_stored2_out & fsm5_out >= 32'd1 & fsm5_out < 32'd4 & fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? tmp_read_data : '0;
  assign t0_in = (fsm2_out == 32'd0 & cond_stored1_out & fsm3_out >= 32'd1 & fsm3_out < 32'd4 & fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? tmp_read_data : '0;
  assign t0_write_en = (fsm2_out == 32'd0 & cond_stored1_out & fsm3_out >= 32'd1 & fsm3_out < 32'd4 & fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? 1'd1 : '0;
  assign tmp_addr0 = (fsm2_out == 32'd0 & cond_stored1_out & fsm3_out >= 32'd1 & fsm3_out < 32'd4 & fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go | fsm6_out == 32'd0 & !tmp_done & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go | fsm2_out == 32'd1 & cond_stored1_out & fsm3_out >= 32'd1 & fsm3_out < 32'd4 & fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go | fsm4_out == 32'd1 & cond_stored2_out & fsm5_out >= 32'd1 & fsm5_out < 32'd4 & fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? i1_out : '0;
  assign tmp_write_data = (fsm6_out == 32'd0 & !tmp_done & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? const6_out : (fsm2_out == 32'd1 & cond_stored1_out & fsm3_out >= 32'd1 & fsm3_out < 32'd4 & fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? add1_out : '0;
  assign tmp_write_en = (fsm6_out == 32'd0 & !tmp_done & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go | fsm2_out == 32'd1 & cond_stored1_out & fsm3_out >= 32'd1 & fsm3_out < 32'd4 & fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? 1'd1 : '0;
  assign x_addr0 = (fsm2_out == 32'd1 & cond_stored1_out & fsm3_out >= 32'd1 & fsm3_out < 32'd4 & fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? j0_out : '0;
  assign y_addr0 = (fsm4_out == 32'd0 & cond_stored2_out & fsm5_out >= 32'd1 & fsm5_out < 32'd4 & fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go | fsm4_out == 32'd1 & cond_stored2_out & fsm5_out >= 32'd1 & fsm5_out < 32'd4 & fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? j1_out : (fsm0_out == 32'd0 & cond_stored0_out & fsm1_out >= 32'd1 & fsm1_out < 32'd3 & fsm7_out == 32'd1 & !(fsm1_out == 32'd1 & !cond_stored0_out) & go) ? i0_out : '0;
  assign y_write_data = (fsm0_out == 32'd0 & cond_stored0_out & fsm1_out >= 32'd1 & fsm1_out < 32'd3 & fsm7_out == 32'd1 & !(fsm1_out == 32'd1 & !cond_stored0_out) & go) ? const2_out : (fsm4_out == 32'd1 & cond_stored2_out & fsm5_out >= 32'd1 & fsm5_out < 32'd4 & fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? add3_out : '0;
  assign y_write_en = (fsm0_out == 32'd0 & cond_stored0_out & fsm1_out >= 32'd1 & fsm1_out < 32'd3 & fsm7_out == 32'd1 & !(fsm1_out == 32'd1 & !cond_stored0_out) & go | fsm4_out == 32'd1 & cond_stored2_out & fsm5_out >= 32'd1 & fsm5_out < 32'd4 & fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? 1'd1 : '0;
  assign y00_in = (fsm4_out == 32'd0 & cond_stored2_out & fsm5_out >= 32'd1 & fsm5_out < 32'd4 & fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? y_read_data : '0;
  assign y00_write_en = (fsm4_out == 32'd0 & cond_stored2_out & fsm5_out >= 32'd1 & fsm5_out < 32'd4 & fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? 1'd1 : '0;
  assign fsm0_in = (fsm0_out != 32'd2 & cond_stored0_out & fsm1_out >= 32'd1 & fsm1_out < 32'd3 & fsm7_out == 32'd1 & !(fsm1_out == 32'd1 & !cond_stored0_out) & go) ? incr0_out : (fsm0_out == 32'd2 & go) ? 32'd0 : '0;
  assign fsm0_write_en = (fsm0_out != 32'd2 & cond_stored0_out & fsm1_out >= 32'd1 & fsm1_out < 32'd3 & fsm7_out == 32'd1 & !(fsm1_out == 32'd1 & !cond_stored0_out) & go | fsm0_out == 32'd2 & go) ? 1'd1 : '0;
  assign incr0_left = (cond_stored0_out & fsm1_out >= 32'd1 & fsm1_out < 32'd3 & fsm7_out == 32'd1 & !(fsm1_out == 32'd1 & !cond_stored0_out) & go) ? 32'd1 : '0;
  assign incr0_right = (cond_stored0_out & fsm1_out >= 32'd1 & fsm1_out < 32'd3 & fsm7_out == 32'd1 & !(fsm1_out == 32'd1 & !cond_stored0_out) & go) ? fsm0_out : '0;
  assign fsm1_in = (fsm1_out != 32'd3 & fsm7_out == 32'd1 & !(fsm1_out == 32'd1 & !cond_stored0_out) & go) ? incr1_out : (fsm1_out == 32'd3 & fsm7_out == 32'd1 & !(fsm1_out == 32'd1 & !cond_stored0_out) & go | fsm1_out == 32'd1 & !cond_stored0_out & go) ? 32'd0 : '0;
  assign fsm1_write_en = (fsm1_out != 32'd3 & fsm7_out == 32'd1 & !(fsm1_out == 32'd1 & !cond_stored0_out) & go | fsm1_out == 32'd3 & fsm7_out == 32'd1 & !(fsm1_out == 32'd1 & !cond_stored0_out) & go | fsm1_out == 32'd1 & !cond_stored0_out & go) ? 1'd1 : '0;
  assign cond_stored0_in = (fsm1_out == 32'd0 & fsm7_out == 32'd1 & !(fsm1_out == 32'd1 & !cond_stored0_out) & go) ? le0_out : '0;
  assign cond_stored0_write_en = (fsm1_out == 32'd0 & fsm7_out == 32'd1 & !(fsm1_out == 32'd1 & !cond_stored0_out) & go) ? 1'd1 : '0;
  assign incr1_left = (fsm7_out == 32'd1 & !(fsm1_out == 32'd1 & !cond_stored0_out) & go) ? fsm1_out : '0;
  assign incr1_right = (fsm7_out == 32'd1 & !(fsm1_out == 32'd1 & !cond_stored0_out) & go) ? 32'd1 : '0;
  assign fsm2_in = (fsm2_out != 32'd3 & cond_stored1_out & fsm3_out >= 32'd1 & fsm3_out < 32'd4 & fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? incr2_out : (fsm2_out == 32'd3 & go) ? 32'd0 : '0;
  assign fsm2_write_en = (fsm2_out != 32'd3 & cond_stored1_out & fsm3_out >= 32'd1 & fsm3_out < 32'd4 & fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go | fsm2_out == 32'd3 & go) ? 1'd1 : '0;
  assign incr2_left = (cond_stored1_out & fsm3_out >= 32'd1 & fsm3_out < 32'd4 & fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? 32'd1 : '0;
  assign incr2_right = (cond_stored1_out & fsm3_out >= 32'd1 & fsm3_out < 32'd4 & fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? fsm2_out : '0;
  assign fsm3_in = (fsm3_out != 32'd4 & fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? incr3_out : (fsm3_out == 32'd4 & fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go | fsm3_out == 32'd1 & !cond_stored1_out & go) ? 32'd0 : '0;
  assign fsm3_write_en = (fsm3_out != 32'd4 & fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go | fsm3_out == 32'd4 & fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go | fsm3_out == 32'd1 & !cond_stored1_out & go) ? 1'd1 : '0;
  assign cond_stored1_in = (fsm3_out == 32'd0 & fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? le2_out : '0;
  assign cond_stored1_write_en = (fsm3_out == 32'd0 & fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? 1'd1 : '0;
  assign incr3_left = (fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? fsm3_out : '0;
  assign incr3_right = (fsm6_out == 32'd2 & !(fsm3_out == 32'd1 & !cond_stored1_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? 32'd1 : '0;
  assign fsm4_in = (fsm4_out != 32'd3 & cond_stored2_out & fsm5_out >= 32'd1 & fsm5_out < 32'd4 & fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? incr4_out : (fsm4_out == 32'd3 & go) ? 32'd0 : '0;
  assign fsm4_write_en = (fsm4_out != 32'd3 & cond_stored2_out & fsm5_out >= 32'd1 & fsm5_out < 32'd4 & fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go | fsm4_out == 32'd3 & go) ? 1'd1 : '0;
  assign incr4_left = (cond_stored2_out & fsm5_out >= 32'd1 & fsm5_out < 32'd4 & fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? 32'd1 : '0;
  assign incr4_right = (cond_stored2_out & fsm5_out >= 32'd1 & fsm5_out < 32'd4 & fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? fsm4_out : '0;
  assign fsm5_in = (fsm5_out != 32'd4 & fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? incr5_out : (fsm5_out == 32'd4 & fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go | fsm5_out == 32'd1 & !cond_stored2_out & go) ? 32'd0 : '0;
  assign fsm5_write_en = (fsm5_out != 32'd4 & fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go | fsm5_out == 32'd4 & fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go | fsm5_out == 32'd1 & !cond_stored2_out & go) ? 1'd1 : '0;
  assign cond_stored2_in = (fsm5_out == 32'd0 & fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? le3_out : '0;
  assign cond_stored2_write_en = (fsm5_out == 32'd0 & fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? 1'd1 : '0;
  assign incr5_left = (fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? fsm5_out : '0;
  assign incr5_right = (fsm6_out == 32'd4 & !(fsm5_out == 32'd1 & !cond_stored2_out) & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? 32'd1 : '0;
  assign fsm6_in = (fsm6_out == 32'd5 & i1_done & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? 32'd6 : (fsm6_out == 32'd4 & fsm5_out == 32'd1 & !cond_stored2_out & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? 32'd5 : (fsm6_out == 32'd3 & j1_done & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? 32'd4 : (fsm6_out == 32'd2 & fsm3_out == 32'd1 & !cond_stored1_out & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? 32'd3 : (fsm6_out == 32'd1 & j0_done & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? 32'd2 : (fsm6_out == 32'd0 & tmp_done & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? 32'd1 : (fsm6_out == 32'd6 & go) ? 32'd0 : '0;
  assign fsm6_write_en = (fsm6_out == 32'd0 & tmp_done & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go | fsm6_out == 32'd1 & j0_done & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go | fsm6_out == 32'd2 & fsm3_out == 32'd1 & !cond_stored1_out & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go | fsm6_out == 32'd3 & j1_done & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go | fsm6_out == 32'd4 & fsm5_out == 32'd1 & !cond_stored2_out & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go | fsm6_out == 32'd5 & i1_done & cond_stored3_out & cond_computed0_out & !(fsm6_out == 32'd6) & fsm7_out == 32'd3 & !(done_reg0_out) & go | fsm6_out == 32'd6 & go) ? 1'd1 : '0;
  assign cond_computed0_in = (cond_stored3_out & cond_computed0_out & fsm6_out == 32'd6 & fsm7_out == 32'd3 & !(done_reg0_out) & go | cond_computed0_out & !cond_stored3_out & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? 1'd0 : (!cond_computed0_out & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? 1'd1 : '0;
  assign cond_computed0_write_en = (!cond_computed0_out & fsm7_out == 32'd3 & !(done_reg0_out) & go | cond_stored3_out & cond_computed0_out & fsm6_out == 32'd6 & fsm7_out == 32'd3 & !(done_reg0_out) & go | cond_computed0_out & !cond_stored3_out & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? 1'd1 : '0;
  assign cond_stored3_in = (!cond_computed0_out & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? le1_out : '0;
  assign cond_stored3_write_en = (!cond_computed0_out & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? 1'd1 : '0;
  assign done_reg0_in = (done_reg0_out & go) ? 1'd0 : (cond_computed0_out & !cond_stored3_out & fsm7_out == 32'd3 & !(done_reg0_out) & go) ? 1'd1 : '0;
  assign done_reg0_write_en = (cond_computed0_out & !cond_stored3_out & fsm7_out == 32'd3 & !(done_reg0_out) & go | done_reg0_out & go) ? 1'd1 : '0;
  assign fsm7_in = (fsm7_out == 32'd3 & done_reg0_out & go) ? 32'd4 : (fsm7_out == 32'd2 & i1_done & go) ? 32'd3 : (fsm7_out == 32'd1 & fsm1_out == 32'd1 & !cond_stored0_out & go) ? 32'd2 : (fsm7_out == 32'd0 & i0_done & go) ? 32'd1 : (fsm7_out == 32'd4 & go) ? 32'd0 : '0;
  assign fsm7_write_en = (fsm7_out == 32'd0 & i0_done & go | fsm7_out == 32'd1 & fsm1_out == 32'd1 & !cond_stored0_out & go | fsm7_out == 32'd2 & i1_done & go | fsm7_out == 32'd3 & done_reg0_out & go | fsm7_out == 32'd4 & go) ? 1'd1 : '0;
endmodule // end main
